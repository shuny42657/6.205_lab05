`default_nettype none
`timescale 1ns / 1ps
module top_level(
	input wire clk,
	input wire btnc,
	input wire[1:0] eth_rxd,
	input wire 

	output logic[15:0] led,

)


`default_nettype wire

